magic
tech sky130A
timestamp 1617838990
<< nmos >>
rect 5 30 20 95
<< ndiff >>
rect -40 80 5 95
rect -40 45 -35 80
rect -15 45 5 80
rect -40 30 5 45
rect 20 80 65 95
rect 20 45 40 80
rect 60 45 65 80
rect 20 30 65 45
<< ndiffc >>
rect -35 45 -15 80
rect 40 45 60 80
<< poly >>
rect 5 95 20 130
rect 5 20 20 30
rect -20 10 20 20
rect -20 -15 -10 10
rect 10 -15 20 10
rect -20 -20 20 -15
<< polycont >>
rect -10 -15 10 10
<< locali >>
rect -90 80 -10 90
rect -90 75 -35 80
rect -90 50 -85 75
rect -65 50 -35 75
rect -90 45 -35 50
rect -15 45 -10 80
rect -90 35 -10 45
rect 35 80 115 90
rect 35 45 40 80
rect 60 75 115 80
rect 60 50 90 75
rect 110 50 115 75
rect 60 45 115 50
rect 35 35 115 45
rect -60 10 20 15
rect -40 -15 -10 10
rect 10 -15 20 10
rect -60 -20 20 -15
<< viali >>
rect -85 50 -65 75
rect 90 50 110 75
rect -60 -15 -40 10
<< metal1 >>
rect -120 75 -55 80
rect -120 50 -85 75
rect -65 50 -55 75
rect -120 45 -55 50
rect 80 75 145 80
rect 80 50 90 75
rect 110 50 145 75
rect 80 45 145 50
rect -95 10 -30 15
rect -95 -15 -60 10
rect -40 -15 -30 10
rect -95 -20 -30 -15
<< labels >>
rlabel metal1 -115 55 -100 70 1 source
rlabel metal1 125 55 140 70 1 drain
rlabel metal1 -85 -10 -70 5 1 gate
<< end >>
