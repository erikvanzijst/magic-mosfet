.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create a resistor between the MOSFET drain and VPWR
R VPWR DRAIN 10k

* create pulse
Vin GATE VGND pulse(0 1.8 100p 10p 10p 500p 1n)
.tran 1p 1n 0

.control
run
set color0 = white
set color1 = black
plot GATE DRAIN
.endc

.end
